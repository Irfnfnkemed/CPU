module alu (
    input wire clk_in,  // system clock signal
    input wire rst_in,  // reset signal
    input wire rdy_in   // ready signal, pause cpu when low
);

endmodule
